----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    03:55:43 04/09/2016 
-- Design Name: 
-- Module Name:    DATA_MEMORY_ADDR_STORAGE - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use ieee.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DATA_MEMORY_ADDR_STORAGE is
PORT(CLK_DEC,CLK_OP,CLK_EX,CLK_WB	 : in STD_LOGIC;
		COUNTER_FOR_WRITING_DATA : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		COUNTER_FOR_OUTPUT_TO_PROCESS: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		COUNTER_FOR_OUTPUT_TO_0_CYCLE_AGO:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		COUNTER_FOR_OUTPUT_TO_1_CYCLE_AGO: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		COUNTER_FOR_OUTPUT_TO_2_CYCLE_AGO: IN STD_LOGIC_VECTOR(2 DOWNTO 0);

		
	
	   DATA_MEMORY_ADDR_IN :in STD_LOGIC_vector(7 downto 0);
		DATA_MEMORY_ADDR_OUT_FOR_PROCESS :out STD_LOGIC_vector(7 downto 0);
		
		DATA_MEMORY_ADDR_OUT_FOR_DATA_0_CYCLE_AGO:out STD_LOGIC_vector(7 downto 0);
		DATA_MEMORY_ADDR_OUT_FOR_DATA_1_CYCLE_AGO:out STD_LOGIC_vector(7 downto 0);
		DATA_MEMORY_ADDR_OUT_FOR_DATA_2_CYCLE_AGO:out STD_LOGIC_vector(7 downto 0)
		


		
		



);
end DATA_MEMORY_ADDR_STORAGE;

architecture Behavioral of DATA_MEMORY_ADDR_STORAGE is
type DATA_MEMORY_ADDR_ARRAY is array (0 to 7) of std_logic_vector(7 downto 0); 
signal DATA_MEMORY_ADDR_SIGNAL : DATA_MEMORY_ADDR_ARRAY:=(0=>"00000000", OTHERS=>"00000000");
signal DATA_MEMORY_ADDR_INTERNAL_SIGNAL_FOR_PROCESS,DATA_MEMORY_ADDR_INTERNAL_SIGNAL_FOR_MEMORY :STD_LOGIC_VECTOR(7 DOWNTO 0);
signal DATA_MEMORY_ADDR_INTERNAL_SIGNAL_FOR_0_CYCLE_AGO,DATA_MEMORY_ADDR_INTERNAL_SIGNAL_FOR_1_CYCLE_AGO,DATA_MEMORY_ADDR_INTERNAL_SIGNAL_FOR_2_CYCLE_AGO :STD_LOGIC_VECTOR(7 DOWNTO 0);
begin

PROCESS(CLK_DEC)
BEGIN
if FALLING_EDGE(CLK_DEC) then
	
		DATA_MEMORY_ADDR_SIGNAL(to_integer(unsigned(COUNTER_FOR_WRITING_DATA)))<=DATA_MEMORY_ADDR_IN;
	
end if;
end process;

with COUNTER_FOR_OUTPUT_TO_PROCESS select
			DATA_MEMORY_ADDR_INTERNAL_SIGNAL_FOR_PROCESS <=
			 DATA_MEMORY_ADDR_SIGNAL(to_integer(unsigned(COUNTER_FOR_OUTPUT_TO_PROCESS)))WHEN "000",
			 DATA_MEMORY_ADDR_SIGNAL(to_integer(unsigned(COUNTER_FOR_OUTPUT_TO_PROCESS)))WHEN OTHERS;
			 
with COUNTER_FOR_OUTPUT_TO_0_CYCLE_AGO select
			DATA_MEMORY_ADDR_INTERNAL_SIGNAL_FOR_0_CYCLE_AGO <=
			 DATA_MEMORY_ADDR_SIGNAL(to_integer(unsigned(COUNTER_FOR_OUTPUT_TO_0_CYCLE_AGO)))WHEN "000",
			 DATA_MEMORY_ADDR_SIGNAL(to_integer(unsigned(COUNTER_FOR_OUTPUT_TO_0_CYCLE_AGO)))WHEN OTHERS;
			 
with COUNTER_FOR_OUTPUT_TO_1_CYCLE_AGO select
			DATA_MEMORY_ADDR_INTERNAL_SIGNAL_FOR_1_CYCLE_AGO <=
			 DATA_MEMORY_ADDR_SIGNAL(to_integer(unsigned(COUNTER_FOR_OUTPUT_TO_1_CYCLE_AGO)))WHEN "000",
			 DATA_MEMORY_ADDR_SIGNAL(to_integer(unsigned(COUNTER_FOR_OUTPUT_TO_1_CYCLE_AGO)))WHEN OTHERS;
			 
with COUNTER_FOR_OUTPUT_TO_2_CYCLE_AGO select
			DATA_MEMORY_ADDR_INTERNAL_SIGNAL_FOR_2_CYCLE_AGO <=
			 DATA_MEMORY_ADDR_SIGNAL(to_integer(unsigned(COUNTER_FOR_OUTPUT_TO_2_CYCLE_AGO)))WHEN "000",
			 DATA_MEMORY_ADDR_SIGNAL(to_integer(unsigned(COUNTER_FOR_OUTPUT_TO_2_CYCLE_AGO)))WHEN OTHERS;


PROCESS(CLK_OP)
BEGIN
if RISING_EDGE(CLK_OP) THEN
		DATA_MEMORY_ADDR_OUT_FOR_DATA_0_CYCLE_AGO<=DATA_MEMORY_ADDR_INTERNAL_SIGNAL_FOR_0_CYCLE_AGO;
		
end if;			 
END PROCESS;

PROCESS(CLK_EX)
BEGIN
if RISING_EDGE(CLK_EX) THEN
		DATA_MEMORY_ADDR_OUT_FOR_DATA_1_CYCLE_AGO<=DATA_MEMORY_ADDR_INTERNAL_SIGNAL_FOR_1_CYCLE_AGO;
		
end if;			 
END PROCESS;


PROCESS(CLK_WB)
BEGIN
if RISING_EDGE(CLK_WB) THEN
		DATA_MEMORY_ADDR_OUT_FOR_DATA_2_CYCLE_AGO<=DATA_MEMORY_ADDR_INTERNAL_SIGNAL_FOR_2_CYCLE_AGO;
		
end if;			 
END PROCESS;

PROCESS(CLK_EX)
BEGIN
if FALLING_EDGE(CLK_EX) THEN
		DATA_MEMORY_ADDR_OUT_FOR_PROCESS<=DATA_MEMORY_ADDR_INTERNAL_SIGNAL_FOR_PROCESS;
end if;			 
END PROCESS;
end Behavioral;

