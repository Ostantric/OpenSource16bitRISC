----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    01:50:41 04/10/2016 
-- Design Name: 
-- Module Name:    DATA_HAZARD_CONTROLLER - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DATA_HAZARD_CONTROLLER is
PORT(

     --SIGNALS_IN
	  CONTROL_IN: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	  control_data_hazard : IN STD_LOGIC;

--CHECK_FLAG:IN STD_LOGIC_VECTOR(3 DOWNTO 0);

--ADDR-------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
     RA_ADDR_2_CYCLE_AGO_IN: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	  RA_ADDR_1_CYCLE_AGO_IN: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	  RA_ADDR_CURRENT_IN,RB_ADDR_CURRENT_IN: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	  DATA_MEMORY_ADDR_1_CYCLE_AGO,DATA_MEMORY_ADDR_2_CYCLE_AGO : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  DATA_MEMORY_ADDR_CURRENT_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  
---DATA_IN-------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	  ALU_RESULT_IN_FOR_1_BYPASS_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	  ALU_RESULT_IN_FOR_2_BYPASS_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	  RA_VALUE_FROM_REG_BANK_IN: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	  RB_VALUE_FROM_REG_BANK_IN: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	  MEM_VALUE_FROM_DATA_MEMORY_IN: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	  EXMEM_VALUE_FROM_EXTERNAL_MEMORY_IN: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	  INSMEM_VALUE_FROM_INSTRUCTION_MEMORY_IN: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	  
--OUT---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	  RA_VALUE_OUT_DATAHAZARD_FIXED : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	  RB_VALUE_OUT_DATAHAZARD_FIXED : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	  MEM_VALUE_OUT_DATAHAZARD_FIXED : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	  EXMEM_VALUE_OUT_DATAHAZARD_FIXED : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	  INSMEM_VALUE_OUT_DATAHAZARD_FIXED: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	  
	  );
end DATA_HAZARD_CONTROLLER;

architecture COMBINATIONAL of DATA_HAZARD_CONTROLLER is
SIGNAL ALU_RESULT_IN_FOR_LOAD_INSTRUCTION,FLAG_CHECK_16BIT : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL RA_VALUE_OUT_DATAHAZARD_FIXED_SIGNAL1,RA_VALUE_OUT_DATAHAZARD_FIXED_SIGNAL2 : STD_LOGIC_VECTOR(15 DOWNTO 0);

begin
--FLAG_CHECK_16BIT<="000000000000" & CHECK_FLAG ;

RA_VALUE_OUT_DATAHAZARD_FIXED<=	ALU_RESULT_IN_FOR_1_BYPASS_IN WHEN RA_ADDR_CURRENT_IN=RA_ADDR_1_CYCLE_AGO_IN ELSE
														ALU_RESULT_IN_FOR_2_BYPASS_IN WHEN RA_ADDR_CURRENT_IN=RA_ADDR_2_CYCLE_AGO_IN ELSE
														RA_VALUE_FROM_REG_BANK_IN;
														
--RA_VALUE_OUT_DATAHAZARD_FIXED_SIGNAL2<=   FLAG_CHECK_16BIT WHEN CONTROL_IN="0010" ELSE
--														X"0000";
--														
--RA_VALUE_OUT_DATAHAZARD_FIXED<= 				RA_VALUE_OUT_DATAHAZARD_FIXED_SIGNAL2 WHEN CONTROL_IN="0010" ELSE
--														RA_VALUE_OUT_DATAHAZARD_FIXED_SIGNAL1;						
					
RB_VALUE_OUT_DATAHAZARD_FIXED<=	ALU_RESULT_IN_FOR_1_BYPASS_IN WHEN RB_ADDR_CURRENT_IN=RA_ADDR_1_CYCLE_AGO_IN ELSE
											ALU_RESULT_IN_FOR_2_BYPASS_IN WHEN RB_ADDR_CURRENT_IN=RA_ADDR_2_CYCLE_AGO_IN ELSE
											RB_VALUE_FROM_REG_BANK_IN;			

ALU_RESULT_IN_FOR_LOAD_INSTRUCTION<=ALU_RESULT_IN_FOR_1_BYPASS_IN	WHEN DATA_MEMORY_ADDR_CURRENT_IN=DATA_MEMORY_ADDR_1_CYCLE_AGO ELSE
												ALU_RESULT_IN_FOR_2_BYPASS_IN WHEN DATA_MEMORY_ADDR_CURRENT_IN=DATA_MEMORY_ADDR_2_CYCLE_AGO ELSE
												MEM_VALUE_FROM_DATA_MEMORY_IN;

											
MEM_VALUE_OUT_DATAHAZARD_FIXED<= ALU_RESULT_IN_FOR_LOAD_INSTRUCTION WHEN control_data_hazard='1' ELSE --LOAD HAZARD FIXED, BUT STILL DIDN'T FIXED THE SPECIAL INSTRUCTION HAZARDS. UPDATE SOON.
											MEM_VALUE_FROM_DATA_MEMORY_IN;



EXMEM_VALUE_OUT_DATAHAZARD_FIXED<=EXMEM_VALUE_FROM_EXTERNAL_MEMORY_IN; -- DATAHAZARD NOT FIXED  YET. JUST NEED ADDTIONAL COMPARING EXMEM ADDRS.

INSMEM_VALUE_OUT_DATAHAZARD_FIXED<=INSMEM_VALUE_FROM_INSTRUCTION_MEMORY_IN;



end COMBINATIONAL;

